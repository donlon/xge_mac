`ifndef XGE_MAC_INCLUDE_SVH
`define XGE_MAC_INCLUDE_SVH

`define transmitData { packetData[7], packetData[6], packetData[5], packetData[4], packetData[3], packetData[2], packetData[1], packetData[0] }

`define receivedData { receivedData [7], receivedData[6], receivedData[5], receivedData[4], receivedData[3], receivedData[2], receivedData[1], receivedData[0] }

`endif